module adder_s_s(
                a,
                b,
                sum
                );
                input [3:0]a;
                input [3:0]b;
                output reg [4:0]sum;
                wire [3:0] internal_sum ;
                assign internal_sum = a + b;
                wire [3:0] a1;   //a�ľ���ֵ
                wire [3:0] b1;   //b�ľ���ֵ
                //һ��һ�����жϾ���ֵ��������ֵ��ȡ0��������ֵ��ȡ1
                //ͬ����ͬ����������λ��0��ֱ�����
                wire [4:0]s_sum;
                assign s_sum = {1'b0,a} + {1'b0,b};
                wire [3:0]c1 ; //���a��b�ķ���
                wire [3:0]c2;
                assign c1 = {1'b0,~a[2:0]};  //���a�ķ���
                assign c2 = {1'b0,~b[2:0]}; //���b�ķ���
                //ȡa��b �ľ���ֵ
                assign a1 = (a[3])  ?  (c1+1) : a[2:0];
                assign b1 = (b[3] ) ?  (c2+1) : b[2:0];
                
                always@(*)begin
                if( (a[3] == 1) &(b[3] == 0)&(a1 >=b1) )
                sum = {1'b1,internal_sum};
                else if( (a[3] == 1) &(b[3] == 0)&(a1 <b1) )
                sum = {1'b0,internal_sum};
                else if((a[3] == 0) & (b[3] == 1) & (a1>=b1) )
                sum = {1'b0,internal_sum};
                else if((a[3] == 0) & (b[3] == 1) & (a1<b1) )
                sum = {1'b1,internal_sum};
                else sum = s_sum;
                end
                
endmodule