module Two_complment #(parameter MIC = 3)(
    in,
    out 
);
        input [MIC-1:0]in;
        output [MIC-1:0]out ;
        //������λ��1����ȡ����һ�������0������ԭֵ
        // //����λ
        // wire sign = in[MIC-1];

        // //����λ
        // wire [MIC-2:0]mag ;
        // assign mag = in[MIC-2:0];
        
        // //���
        // assign out = sign ? {1'b1,~mag+1} : in;
        
        
        //�򻯰��
assign out = in[MIC-1] ? {1'b1,{~in[MIC-2:0]+1}} : in;

endmodule 